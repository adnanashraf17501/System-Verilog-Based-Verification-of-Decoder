`ifndef base_pkt
`define base_pkt
class base_pkt;
           rand bit [3:0]x;
	       bit [15:0]y;
	bit en;
endclass 
`endif
